--create 4 bit adder

--test bench definition
--Port( X: in STD_logic
--      B
--      ci<= test(8)
    wat9f f0r
